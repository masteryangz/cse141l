111111111 //mem[64] = 64
110000111 //r0 = 64
110001111 //r1 = 64
111010111 //max(mem[64]) = 0
001000001 //r0 = 32
001000001 //r0 = 16
010111110 //r7 = 65
111000111 //min(mem[65]) = 16
010111110 //r7 = 66
111010111 //mem[66] = 0
010111110 //r7 = 67
111001111 //mem[67] = 64
010111110 //r7 = 68
010111110 //r7 = 69
111101111 //mem[69] = -1
010111110 //r7 = 70
111110111 //mem[70] = 1
110111111 //r7 = 64
110000111 //r0 = 0
110001111 //r1 = 0
110011111 //r3 = 0
010011010 //load r3 with r2(i)
100011101 //r3 = ~r2
010011110 //r3 = -r2
010111101 //r7 = len(n)-1
010111101 //r7 = len(n)-2
010011111 //r3 = len(n)-2-i
010111110 //r7 = len(n)-1
010111110 //r7 = len(n)
101011110 //for i in range(len(n)-1)
010111110 //r7 = len(n)+1
010111110 //r7 = len(n)+2
110011111 //r3 = 0
010011110 //r3 = 1
010011110 //r3 = 2
010011010 //r3(j) = r2(i)+2
110100111 //r4 = 0
010100011 //load r4 with r3(j)
100100101 //r4 = ~r3
010100110 //r4 = -r3
010111101 //r7 = len(n)+1
010111101 //r7 = len(n)
010111101 //r7 = len(n)-1
010100111 //r4 = len(n)-1-j
010111110 //r7 = len(n)
101100100 //for j in range(i+1, len(n))
110100010 //load mem[i] into r4
110000011 //load mem[j] into r0
100100101 //r4 = ~r4
010100110 //r4 = r4+1(-mem[j])
010000100 //r0(setBits) = r0(mem[i])+r4(-mem[j])
011000010 //if r0(setBits)<0
100000101 //r0 = ~r0
010000110 //r0 = r0+1(-setBits)
010011110 //j+=1
010011110 //j+=1
101101101 //jump back to j for loop
010010110 //i+=1
010010110 //i+=1
101101111 //jump back to i for loop
