000000110 //line1
010110100 //line2
