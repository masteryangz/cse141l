111111111 //mem[64] = 64
110000111 //r0 = 64
110001111 //r1 = 64
111010111 //max(mem[64]) = 0
001000001 //r0 = 32
001000001 //r0 = 16
010111110 //r7 = 65
111000111 //min(mem[65]) = 16
010111110 //r7 = 66
111010111 //mem[66] = 0
010111110 //r7 = 67
111001111 //mem[67] = 64
010111110 //r7 = 68
111101111 //mem[68] = -1
010111110 //r7 = 69
111110111 //mem[69] = 1
010111110 //r7 = 68
010111110 //r7 = 67
010111110 //r7 = 66
010111110 //r7 = 65
010111110 //r7 = 64
110000111 //r0 = mem[64](0)
110001111 //r1 = mem[64](0)
110011111 //r3 = mem[64](0)