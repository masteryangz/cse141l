010000001 //line1
000011010 //line2
001000101 //line3
011000011 //line4
100111110 //line5
101011101 //line6
110001000 //line7
111000001 //line8
111000001 //line9
